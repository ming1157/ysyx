
package arb_pkg;

//arbiter package
  class arb_trans;
    // ... ignored
  endclass

  class arb_driver;
    // ... ignored
  endclass

  class arb_generator;
    // ... ignored
  endclass

  class arb_monitor;
    // ... ignored
  endclass

  class arb_agent;
    // ... ignored
  endclass
endpackage

